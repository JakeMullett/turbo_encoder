module read_fsm();

endmodule
